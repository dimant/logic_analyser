   event t_fail;
   
   always @(t_fail)
     $display("FAIL");   
